library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
	port(
		addr : in std_logic_vector(8 downto 0);
		data : out std_logic_vector(16 downto 0)
		);
	end ROM;

architecture LUT of ROM is
begin
	process(addr)
	begin
		case addr is
			when "000000000" => data <= "10000010100001110";
			when "000000001" => data <= "10111111100001110";
			when "000000010" => data <= "10111101000000110";
			when "000000011" => data <= "10111111100001100";
			when "000000100" => data <= "00001010000011101";
			when "000000101" => data <= "10111101000000010";
			when "000000110" => data <= "10111111100001101";
			when "000000111" => data <= "00001010000011101";
			when "000001000" => data <= "10111101000000011";
			when "000001001" => data <= "10111111100001110";
			when "000001010" => data <= "00001010000011101";
			when "000001011" => data <= "10111101000000100";
			when "000001100" => data <= "00001010001000111";
			when "000001101" => data <= "10000010100001100";
			when "000001110" => data <= "11111100100001010";
			when "000001111" => data <= "10100000100001100";
			when "000010000" => data <= "00010010000000000";
			when "000010001" => data <= "10110010000001100";
			when "000010010" => data <= "10000010100001101";
			when "000010011" => data <= "11111100100001010";
			when "000010100" => data <= "10100000100001101";
			when "000010101" => data <= "00010010000000000";
			when "000010110" => data <= "10110010000001101";
			when "000010111" => data <= "10000010100001110";
			when "000011000" => data <= "11111100100001010";
			when "000011001" => data <= "10100000100001110";
			when "000011010" => data <= "00010010000000000";
			when "000011011" => data <= "10110010000001110";
			when "000011100" => data <= "00010010000000000";
			when "000011101" => data <= "10111101000001011";
			when "000011110" => data <= "11111100100000000";
			when "000011111" => data <= "10100001000001011";
			when "000100000" => data <= "00010010000111101";
			when "000100001" => data <= "11111100100000001";
			when "000100010" => data <= "10100001000001011";
			when "000100011" => data <= "00010010000111110";
			when "000100100" => data <= "11111100100000010";
			when "000100101" => data <= "10100001000001011";
			when "000100110" => data <= "00010010000111111";
			when "000100111" => data <= "11111100100000011";
			when "000101000" => data <= "10100001000001011";
			when "000101001" => data <= "00010010001000000";
			when "000101010" => data <= "11111100100000100";
			when "000101011" => data <= "10100001000001011";
			when "000101100" => data <= "00010010001000001";
			when "000101101" => data <= "11111100100000101";
			when "000101110" => data <= "10100001000001011";
			when "000101111" => data <= "00010010001000010";
			when "000110000" => data <= "11111100100000110";
			when "000110001" => data <= "10100001000001011";
			when "000110010" => data <= "00010010001000011";
			when "000110011" => data <= "11111100100000111";
			when "000110100" => data <= "10100001000001011";
			when "000110101" => data <= "00010010001000100";
			when "000110110" => data <= "11111100100001000";
			when "000110111" => data <= "10100001000001011";
			when "000111000" => data <= "00010010001000101";
			when "000111001" => data <= "11111100100001001";
			when "000111010" => data <= "10100001000001011";
			when "000111011" => data <= "00010010001000110";
			when "000111100" => data <= "00110000000000000";
			when "000111101" => data <= "00101010000000001";
			when "000111110" => data <= "00101010001001111";
			when "000111111" => data <= "00101010000010010";
			when "001000000" => data <= "00101010000000110";
			when "001000001" => data <= "00101010001001100";
			when "001000010" => data <= "00101010000100100";
			when "001000011" => data <= "00101010000100000";
			when "001000100" => data <= "00101010000001111";
			when "001000101" => data <= "00101010000000000";
			when "001000110" => data <= "00101010000001100";
			when "001000111" => data <= "10000111000001000";
			when "001001000" => data <= "00010010001000111";
			when "001001001" => data <= "10000111000001001";
			when "001001010" => data <= "00010010001000111";
			when "001001011" => data <= "10000111000001010";
			when "001001100" => data <= "00010010001000111";
			when "001001101" => data <= "00110000000000000";
			when others => data <= "00000000000000000";
		end case;
	end process;
end LUT;
